module Adder(input logic [31:0] input0,input1, output logic [31:0] out);
assign out = input0 + input1;
endmodule